module clock_divider